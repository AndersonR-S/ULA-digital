library verilog;
use verilog.vl_types.all;
entity MRB_vlg_vec_tst is
end MRB_vlg_vec_tst;
