library verilog;
use verilog.vl_types.all;
entity registradores_32bits_vlg_vec_tst is
end registradores_32bits_vlg_vec_tst;
