library verilog;
use verilog.vl_types.all;
entity memoria_RAM_vlg_vec_tst is
end memoria_RAM_vlg_vec_tst;
