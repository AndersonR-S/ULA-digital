library verilog;
use verilog.vl_types.all;
entity ULA_32_vlg_vec_tst is
end ULA_32_vlg_vec_tst;
